LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY ContadorBCD IS
	PORT(
		MX_CNT, MI_CNT: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		STP_CNT: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		UPDW_CNT, CK_CNT, CLR_CNT: IN STD_LOGIC;
		Q_CNT: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
		LED_CNT: OUT STD_LOGIC
	);
END ContadorBCD;

ARCHITECTURE contador OF ContadorBCD IS
	
	COMPONENT RegistradorAcumulador IS
		PORT(
			A_RA: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			CK_RA, CLR_RA: IN STD_LOGIC;
			Q_RA: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT SomadorBCD IS
		PORT(
			A_BCD, B_BCD: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			CI_BCD: IN STD_LOGIC;
			S_BCD: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			CO_BCD: OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT Somador4Bits IS
    PORT(
        A_S4B, B_S4B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        CI_S4B: IN STD_LOGIC;
        S_S4B: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
        CO_S4B: OUT STD_LOGIC
    );
	END COMPONENT;
	
	COMPONENT Subtrator IS
		PORT(
			A_SUC, B_SUC: IN STD_LOGIC_VECTOR (3 DOWNTO 0); 
			TI_SUC: IN STD_LOGIC;
			S_SUC: OUT STD_LOGIC_VECTOR (3 DOWNTO 0) ;
			TO_SUC: OUT STD_LOGIC
		);
	END COMPONENT;	
	
	COMPONENT COMPARADOR is

		port(A_mx,B_mn,S_C: in std_logic_vector(11 downto 0);updw : std_logic;igual: out std_logic);

	end COMPONENT;

	SIGNAL Q_REG, D_REG, D_SUM, D_SUB: STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
	SIGNAL CO_CNT, TO_CNT: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL UPDW_VEC: STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
	SIGNAL COMP_UN, COMP_DE: STD_LOGIC;
	SIGNAL Q_CORR_UN, Q_CORR_DE, Q_CORR_CE, V_CORR, STP_CORR: STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL COMP_VEC_DE: STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL COUT_T, EN_STP: STD_LOGIC;
	SIGNAL STP_FINAL, EN_STP_VEC: STD_LOGIC_VECTOR (3 DOWNTO 0);
	
BEGIN 
R0: RegistradorAcumulador PORT MAP(D_REG, CK_CNT, CLR_CNT, Q_REG);

COMP: COMPARADOR PORT MAP(MX_CNT, MI_CNT, Q_REG, UPDW_CNT, EN_STP);
LED_CNT <= EN_STP;
EN_STP_VEC <= (OTHERS => EN_STP);
STP_FINAL <= (STP_CNT AND NOT EN_STP_VEC) OR ("0000" AND EN_STP_VEC);

C0: SomadorBCD PORT MAP(Q_REG(3 DOWNTO 0), STP_FINAL, '0', D_SUM(3 DOWNTO 0), CO_CNT(0));
C1: SomadorBCD PORT MAP(Q_REG(7 DOWNTO 4), "0000", CO_CNT(0), D_SUM(7 DOWNTO 4), CO_CNT(1));
C2: SomadorBCD PORT MAP(Q_REG(11 DOWNTO 8), "0000", CO_CNT(1), D_SUM(11 DOWNTO 8), CO_CNT(2));

COMP_UN <=  (not(Q_REG(3)) and STP_FINAL(3)) or 
((Q_REG(3) xnor STP_FINAL(3)) and not(Q_REG(2)) and STP_FINAL(2) ) or 
((Q_REG(3) xnor STP_FINAL(3)) and (Q_REG(2) xnor STP_FINAL(2)) and  not(Q_REG(1)) and STP_FINAL(1)) or 
((Q_REG(3) xnor STP_FINAL(3)) and (Q_REG(2) xnor STP_FINAL(2)) and  
(Q_REG(1) xnor STP_FINAL(1)) and  not(Q_REG(0)) and STP_FINAL(0));

V_CORR(1) <= COMP_UN;
V_CORR(3) <= COMP_UN;

SUM_CORR: Somador4Bits PORT MAP(Q_REG(3 DOWNTO 0), V_CORR, '0', Q_CORR_UN, COUT_T);

SUB0: Subtrator PORT MAP(Q_CORR_UN, STP_FINAL, '0', D_SUB(3 DOWNTO 0), TO_CNT(0));

STP_CORR(0) <= ('0' AND NOT(COMP_UN)) OR ('1' AND COMP_UN);
COMP_DE <= NOT(Q_REG(7)) AND NOT(Q_REG(6)) AND NOT(Q_REG(5)) AND NOT(Q_REG(4)) AND 
				NOT(STP_CORR(3)) AND NOT(STP_CORR(2)) AND NOT(STP_CORR(1)) AND STP_CORR(0);
COMP_VEC_DE <= (OTHERS => COMP_DE);
Q_CORR_DE <= (Q_REG(7 DOWNTO 4) AND NOT(COMP_VEC_DE)) OR ("1010" AND COMP_VEC_DE);

SUB1: Subtrator PORT MAP(Q_CORR_DE, STP_CORR, '0', D_SUB(7 DOWNTO 4), TO_CNT(1));
SUB2: Subtrator PORT MAP(Q_REG(11 DOWNTO 8), ("0000" AND NOT(COMP_VEC_DE)) OR ("0001" AND COMP_VEC_DE), '0', D_SUB(11 DOWNTO 8), TO_CNT(2));

UPDW_VEC <= (OTHERS => UPDW_CNT);
D_REG <= (D_SUB AND NOT UPDW_VEC) OR (D_SUM AND UPDW_VEC);
Q_CNT <= D_REG;

END contador;